module EX_to_WB
  (


  );




endmodule