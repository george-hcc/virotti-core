package ctrl_typedefs;

typedef enum
  {
    OP_NO_OP,
    OP_COMP,
    OP_COMP_IMM,
    OP_STORE,
    OP_LOAD,
    OP_BRANCH,
    OP_JALR,
    OP_JAL,
    OP_AUIPC,
    OP_LUI,
  } decoded_opcode;

typedef enum
  {
    INSTR_NO_OP,
    INSTR_ADD,
    INSTR_SUB,
    INSTR_SLL,
    INSTR_SRL,
    INSTR_SRA,
    INSTR_AND,
    INSTR_OR,
    INSTR_XOR,
    INSTR_SLT,
    INSTR_SLTU,
    INSTR_ADDI,
    INSTR_SLLI,
    INSTR_SRLI,
    INSTR_SRAI,
    INSTR_ANDI,
    INSTR_ORI,
    INSTR_XORI,
    INSTR_SLTI,
    INSTR_SLTIU,
    INSTR_LUI,
    INSTR_AUIPC,
    INSTR_LB,
    INSTR_LBU,
    INSTR_LH,
    INSTR_LHU,
    INSTR_LW,
    INSTR_SB,
    INSTR_SH,
    INSTR_SW,
    INSTR_FENCE,
    INSTR_FENCEI,
    INSTR_BEQ,
    INSTR_BNE,
    INSTR_BLT,
    INSTR_BLTU,
    INSTR_BGE,
    INSTR_BGEU,
    INSTR_JAL,
    INSTR_JALR,
    INSTR_MUL,
    INSTR_MULH,
    INSTR_MULHSU,
    INSTR_MULHU,
    INSTR_DIV,
    INSTR_DIVU,
    INSTR_REM,
    INSTR_REMU,
    INSTR_BAD_INSTR
  } decoded_instr;

endpackage