module ID_EX_FF
  (

  );





endmodule