module ID_to_EX
  (

  );





endmodule