module IF_to_ID
  (


  );



endmodule